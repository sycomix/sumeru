../../libsrc/alt_ram.vhd